* EESchema Netlist Version 1.1 (Spice format) creation date: 12/03/2015 17:06:55

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
P1_STM1  GNDPWR GNDPWR VDD VDD GNDPWR ? ? ? ? ? ? PA0 PA3 PA2 PA5 ? ? ? ? ? PB1 PB0 GNDPWR ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? GNDPWR GNDPWR CONN_02X25		
P2_STM1  GNDPWR GNDPWR +5V +5V +3V3 +3V3 ? ? ? ? ? ? ? ? ? ? ? ? ? PB9 ? VDD ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? PC6 ? GNDPWR GNDPWR CONN_02X25		
P3_SERVO1  GNDPWR +5C PA3 CONN_01X03		
P4_SERVO1  GNDPWR +5C PA5 CONN_01X03		
P6_SERVO1  GNDPWR +5C PB0 CONN_01X03		
P5_SERVO1  GNDPWR +5C PB1 CONN_01X03		
D2  Net-_D2-Pad1_ ? DIODE		
P1_POL1  ? ? CONN_01X02		
P2_POL1  ? ? CONN_01X02		
P3_POL1  ? ? CONN_01X02		
P4-_POL1  ? ? CONN_01X02		
D3  Net-_D3-Pad1_ ? DIODE		
D4  Net-_D4-Pad1_ ? DIODE		
D5  Net-_D5-Pad1_ ? DIODE		
D1  Net-_D1-Pad1_ ? DIODE		
P2_SERVO1  GNDPWR +5C PA2 CONN_01X03		
P1_SERVO1  GNDPWR +5C PA0 CONN_01X03		
P6_POL1  ? ? CONN_01X02		
P5_POL1  ? ? CONN_01X02		
R2  Net-_D2-Pad1_ ? R		
R3  ? Net-_D3-Pad1_ R		
R4  ? Net-_D4-Pad1_ R		
R5  ? Net-_D5-Pad1_ R		
R1  ? Net-_D1-Pad1_ R		
P7_SERVO1  GNDPWR +5C PC6 CONN_01X03		
P8_SERVO1  GNDPWR +5C PB9 CONN_01X03		
P7_POL1  ? ? CONN_01X02		
P8_POL1  ? ? CONN_01X02		

.end
